    ����          Assembly-CSharp   �System.Collections.Generic.List`1[[Input_text+Tabl_rec, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  Input_text+Tabl_rec[]   	                   Input_text+Tabl_rec      Input_text+Tabl_rec   namescore       ыыы            ффф         
    	      
     