    ����          Assembly-CSharp   Next_level+Saver   level       