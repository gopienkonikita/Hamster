    ����          Assembly-CSharp   Menu_pause+Saver   lvlxyzhealthcoins
bonus_jump             ,��f��              